module Q2_2
(
	input a, b,
	output s, c
);

//assignments...

assign s = a ^ b;

assign c = a & b;

endmodule